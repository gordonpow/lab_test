library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PWM_Generator is
    Port (
        clk     : in  STD_LOGIC;          -- �t�ή���
        reset   : in  STD_LOGIC;          -- �D�P�B���]
        input_n : in  unsigned(3 downto 0); -- ��J�� (1, 2, 3...)
        pwm_out : out STD_LOGIC           -- PWM ��X�H��
    );
end PWM_Generator;

architecture Behavioral of PWM_Generator is
    -- ���]�p�ƾ��q 0 �� 9 (�@ 10 �Ӷ��h)
    signal counter : unsigned(3 downto 0) := (others => '0');
begin
    process(clk, reset)
    begin
        if reset = '1' then
            counter <= (others => '0');
            pwm_out <= '0';
        elsif rising_edge(clk) then
            -- �p�ƾ��b 0-9 �����`��
            if counter >= 9 then
                counter <= (others => '0');
            else
                counter <= counter + 1;
            end if;

            -- ����޿�G��p�ƾ��p���J�ȮɡA��X���q��
            -- �Ҧp input_n = 1�A�h�� counter = 0 �ɿ�X '1' (�e 1/10 = 10%)
            if counter < input_n then
                pwm_out <= '1';
            else
                pwm_out <= '0';
            end if;
        end if;
    end process;
end Behavioral;