library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_Random_Gen is
-- Testbench ���ݭn Port
end tb_Random_Gen;

architecture sim of tb_Random_Gen is
    -- �ŧi�P����ۦP���T��
    signal clk      : std_logic := '0';
    signal reset    : std_logic := '0';
    signal input_en : std_logic := '0';
    signal rand_out : std_logic_vector(1 downto 0);

    -- �w�q�����g�� (10ns = 100MHz)
    constant clk_period : time := 10 ns;

begin
    -- ��ҤƳQ������ (UUT)
    uut: entity work.Random_Gen_0to3
        port map (
            clk      => clk,
            reset    => reset,
            input_en => input_en,
            rand_out => rand_out
        );

    -- �i�קﳡ���j�L���`�����������͹L�{
    clk_process : process
    begin
        clk <= '0';
        wait for clk_period / 2;
        clk <= '1';
        wait for clk_period / 2;
        -- �o�̤��ݭn loop�Aprocess �������槹�N�|�q�Y�}�l�A�F���L�� CLK
    end process;

    -- ��E�L�{ (Stimulus process)
    stim_proc: process
    begin		
        -- 1. �t�έ��m
        reset <= '0';
        wait for 22 ns; -- �y�L�����A�׶}�W�ɪu�H�T�O�T��í�w
        reset <= '1';
        wait for clk_period;

        -- 2. �]�w��J�� 1�A�}�l�ͦ��H����
        input_en <= '1';
        
        -- ����@�q�ɶ��H���ͳs���H����
        -- �Y�n�b�������ݨ쵲�G�A�Ф�ʳ]�w��������ɶ� (�p run 1us)
        wait for clk_period * 10; 

        -- 3. ����ͦ�
        input_en <= '0';
        
        -- �����N�|�b�o�̫��򱾰_�A�� clk_process �|�b�I���@������
        wait; 
    end process;

end sim;