library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Random_Gen_0to3 is
    Port (
        clk      : in  STD_LOGIC;
        reset    : in  STD_LOGIC;
        input_en : in  STD_LOGIC;
        rand_out : out STD_LOGIC_VECTOR(1 downto 0) -- �D�حn�D��X q[0]�A�o�̨���찵 0-3
    );
end Random_Gen_0to3;

architecture Behavioral of Random_Gen_0to3 is
    -- �ھڹϤ��D�ءG��l�Ȭ� 11110
    signal q : std_logic_vector(4 downto 0) := "11110"; 
begin
    process(clk, reset)
    begin
        if reset = '0' then
            q <= "11110"; -- �D�حn�D�� Reset ��
        elsif falling_edge(clk) then
            if input_en = '1' then
                q(4) <= q(0) xor '0';      -- �̥��䪺 XOR (�� 0)
                q(3) <= q(4);              -- ��������
                q(2) <= q(3) xor q(0);     -- ������ XOR (q[3] xor q[0])
                q(1) <= q(2);              -- ��������
                q(0) <= q(1);              -- ��������
            end if;
        end if;
    end process;

    -- ��X�M�g�G�D�ػ���X�b q[0]�A�Y�n�ͦ� 0-3�A�ڭ̨� q(1 downto 0)
    rand_out <= q(1 downto 0);
end Behavioral;