library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity PWM_Generator_tb is
-- Testbench ���ݭn Port
end PWM_Generator_tb;

architecture sim of PWM_Generator_tb is
    -- �ŧi�P����ۦP���T��
    signal clk     : std_logic := '0';
    signal reset   : std_logic := '0';
    signal input_n : unsigned(3 downto 0) := (others => '0');
    signal pwm_out : std_logic;

    -- �w�q�����g�� (�Ҧp 100MHz = 10ns)
    constant clk_period : time := 10 ns;

begin
    -- ��ҤƳQ������ (UUT)
    uut: entity work.PWM_Generator
        port map (
            clk     => clk,
            reset   => reset,
            input_n => input_n,
            pwm_out => pwm_out
        );

    -- �������͹L�{
    clk_process : process
    begin
        while now < 1000 ns loop  -- �`�@���� 1000ns
            clk <= '0';
            wait for clk_period / 2;
            clk <= '1';
            wait for clk_period / 2;
        end loop;
        wait;
    end process;

    -- ��E�L�{ (Stimulus process)
    stim_proc: process
    begin		
        -- 1. ��l�ƻP���]
        reset <= '1';
        wait for 20 ns;
        reset <= '0';

        -- 2. ���� 10% �e�Ť� (Input = 1)
        input_n <= "0001";
        wait for 150 ns;

        -- 3. ���� 20% �e�Ť� (Input = 2)
        input_n <= "0010";
        wait for 150 ns;

        -- 4. ���� 50% �e�Ť� (Input = 5)
        input_n <= "0101";
        wait for 150 ns;

        -- �������
        wait;
    end process;

end sim;