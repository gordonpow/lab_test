library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity traffic_light_fsm_tb is
-- Testbench ���ݭn�� (Ports)
end traffic_light_fsm_tb;

architecture sim of traffic_light_fsm_tb is

    -- �ŧi�ݴ����� (UUT)
    component traffic_light_fsm
        Port ( 
            clk   : in  STD_LOGIC;
            rst_n : in  STD_LOGIC;
            light : out STD_LOGIC_VECTOR (2 downto 0)
        );
    end component;

    -- �����T���ŧi
    signal clk   : STD_LOGIC := '0';
    signal rst_n : STD_LOGIC := '0';
    signal light : STD_LOGIC_VECTOR (2 downto 0);

    -- �ɯ߶g���w�q (10ns = 100MHz)
    constant clk_period : time := 10 ns;

begin

    -- ����ƫݴ����� (Unit Under Test)
    uut: traffic_light_fsm Port map (
          clk   => clk,
          rst_n => rst_n,
          light => light
        );

    -- �ɯ߲��͵{��
    clk_process : process
    begin
        while now < 500 ns loop -- �������� 500ns �ᰱ��
            clk <= '0';
            wait for clk_period/2;
            clk <= '1';
            wait for clk_period/2;
        end loop;
        wait;
    end process;

    -- ���տE�y�{�� (Stimulus Process)
    stim_proc: process
    begin		
        -- ��l���A�G���m�t��
        rst_n <= '0';
        wait for 20 ns;	
        
        rst_n <= '1'; -- ���񭫸m�A�}�l�B�@
        
        -- �[��i���ഫ
        -- ��O������ 80ns (8 clks * 10ns)
        -- ���O������ 20ns (2 clks * 10ns)
        -- ���O������ 100ns (10 clks * 10ns)
        
        wait;
    end process;

end sim;